`timescale 1 ps / 1 ps

module design_1_wrapper
   (y_0);
  output y_0;

  wire y_0;

  design_1 design_1_i
       (.y_0(y_0));
endmodule
